// mem types
parameter int PROC_MEM_TYPE_RAM = 0;
parameter int PROC_MEM_TYPE_REG = 1;
parameter int PROC_MEM_TYPE_STK = 2;
parameter int PROC_MEM_TYPE_COUNT = 3;

parameter int DEBUG_MEM_TYPE_RAM = 0;
parameter int DEBUG_MEM_TYPE_VRAM = 1;
parameter int DEBUG_MEM_TYPE_REG = 2;
parameter int DEBUG_MEM_TYPE_STK = 3;
parameter int DEBUG_MEM_TYPE_COUNT = 4;
