// mem types
parameter int PROC_MEM_TYPE_RAM = 0;
parameter int PROC_MEM_TYPE_REG = 1;
parameter int PROC_MEM_TYPE_STK = 2;
parameter int PROC_MEM_TYPE_COUNT = 3;

parameter int DEBUG_MEM_TYPE_RAM = 0;
parameter int DEBUG_MEM_TYPE_VRAM = 1;
parameter int DEBUG_MEM_TYPE_REG = 2;
parameter int DEBUG_MEM_TYPE_STK = 3;
parameter int DEBUG_MEM_TYPE_COUNT = 4;

parameter int VIDEO_MEM_TYPE_RAM = 0;
parameter int VIDEO_MEM_TYPE_VRAM = 1;
parameter int VIDEO_MEM_TYPE_COUNT = 2;

parameter int REG_V0 = 0;
parameter int REG_V1 = 1;
parameter int REG_V2 = 2;
parameter int REG_V3 = 3;
parameter int REG_V4 = 4;
parameter int REG_V5 = 5;
parameter int REG_V6 = 6;
parameter int REG_V7 = 7;
parameter int REG_V8 = 8;
parameter int REG_V9 = 9;
parameter int REG_VA = 10;
parameter int REG_VB = 11;
parameter int REG_VC = 12;
parameter int REG_VD = 13;
parameter int REG_VE = 14;
parameter int REG_VF = 15;
parameter int REG_I  = 16;
parameter int REG_PC = 18;
parameter int REG_SP = 20;
parameter int REG_DT = 21;
parameter int REG_ST = 22;
