// mem types
parameter int PROC_MEM_TYPE_RAM = 0;
parameter int PROC_MEM_TYPE_REG = 1;
parameter int PROC_MEM_TYPE_STK = 2;
